import uvm_pkg::*;
`include "uvm_macros.svh"

import svt_uvm_pkg::*;

//`default_nettype none
//
//`include "svt_i2c.uvm.pkg"
//`include "i2c_mstr1_i2c_system_configuration.sv"
//`include "i2c_slv1_i2c_system_configuration.sv"
//`include "tb_env.sv"
