
`include "i2c_master_seq_item.sv"
`include "i2c_slave_seq_item.sv"
`include "i2c_sequence_lib.sv"
`include "base_sequence.sv"
`include "basic_bmc_side_rw_seq.sv"

