`include "base_test.sv"
`include "basic_bmc_side_rw_test.svh"
